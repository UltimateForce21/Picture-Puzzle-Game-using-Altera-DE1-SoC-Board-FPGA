/******************************************************************************
 *                                                                            *
 * Module:       Hexadecimal_To_Seven_Segment                                 *
 * Description:                                                               *
 *      This module converts hexadecimal numbers for seven segment displays.  *
 *                                                                            *
 ******************************************************************************/

module Hexadecimal_To_Seven_Segment (
	// Inputs
	hex_number,

	// Bidirectional

	// Outputs
	seven_seg_display
);

/*****************************************************************************
 *                           Parameter Declarations                          *
 *****************************************************************************/


/*****************************************************************************
 *                             Port Declarations                             *
 *****************************************************************************/
// Inputs
input		[2:0]	hex_number;

// Bidirectional

// Outputs
output		[6:0]	seven_seg_display;

/*****************************************************************************
 *                 Internal Wires and Registers Declarations                 *
 *****************************************************************************/
// Internal Wires

// Internal Registers

// State Machine Registers

/*****************************************************************************
 *                         Finite State Machine(s)                           *
 *****************************************************************************/


/*****************************************************************************
 *                             Sequential Logic                              *
 *****************************************************************************/


/*****************************************************************************
 *                            Combinational Logic                            *
 *****************************************************************************/

assign seven_seg_display =
		({7{(hex_number == 3'd0)}} & 7'b1000000) |
		({7{(hex_number == 3'd1)}} & 7'b1111001) |
		({7{(hex_number == 3'd2)}} & 7'b0100100) |
		({7{(hex_number == 3'd3)}} & 7'b0110000) |
		({7{(hex_number == 3'd4)}} & 7'b0011001) |
		({7{(hex_number == 3'd5)}} & 7'b1001110); 

/*****************************************************************************
 *                              Internal Modules                             *
 *****************************************************************************/


endmodule


//assign seven_seg_display =
//		({7{(hex_number == 3'd0)}} & 7'b1000000) |
//		({7{(hex_number == 3'd1)}} & 7'b1111001) |
//		({7{(hex_number == 3'd2)}} & 7'b0100100) |
//		({7{(hex_number == 3'd3)}} & 7'b0110000) |
//		({7{(hex_number == 3'd4)}} & 7'b0011001) |
//		({7{(hex_number == 3'd5)}} & 7'b0010010) |
//		({7{(hex_number == 4'h6)}} & 7'b0000010) |
//		({7{(hex_number == 4'h7)}} & 7'b1111000) |
//		({7{(hex_number == 4'h8)}} & 7'b0000000) |
//		({7{(hex_number == 4'h9)}} & 7'b0010000) |
//		({7{(hex_number == 4'hA)}} & 7'b0001000) |
//		({7{(hex_number == 4'hB)}} & 7'b0000011) |
//		({7{(hex_number == 4'hC)}} & 7'b1000110) |
//		({7{(hex_number == 4'hD)}} & 7'b0100001) |
//		({7{(hex_number == 4'hE)}} & 7'b0000110) |
//		({7{(hex_number == 4'hF)}} & 7'b0001110); 

